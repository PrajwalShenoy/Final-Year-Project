`timescale 1ns / 1ps

module andg16_tb();
reg [15:0]x,y;
wire [15:0]out;
and16 and1(out,x,y);
initial begin
x = 16'b0000000000000000; y = 16'b0000000000000000;#5
x = 16'b0000000000000000; y = 16'b0000000000000001;#5
x = 16'b0000000000000011; y = 16'b0000000000000001;#5
x = 16'b0000000000001111; y = 16'b1111100000001111;#5
$finish;
end
endmodule